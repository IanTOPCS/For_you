library verilog;
use verilog.vl_types.all;
entity tb_accumulator_top is
end tb_accumulator_top;
