`timescale 1ns/100ps
module Program_Rom(
	input	logic [31:0] Rom_addr,
	output	logic [31:0] Rom_data
);    
  
    always_comb begin
        case (Rom_addr)
			32'h0  : Rom_data = 32'h00100093;	//addi	x1, x0, 1	
			32'h4  : Rom_data = 32'h00200113;	//addi	x2, x0, 2	
			32'h8  : Rom_data = 32'hffd00193;	//addi	x3, x0, -3
			32'hc  : Rom_data = 32'h0060a213;	//slti	x4, x1, 6    
			32'h10 : Rom_data = 32'h0060b293;	//sltiu	x5, x1, 6   
			32'h14 : Rom_data = 32'h7ff0f313;	//andi  x6, x1, 2047
			32'h18 : Rom_data = 32'h7ff16393;	//ori   x7, x2, 2047
			32'h1c : Rom_data = 32'h7ff1c413;	//xori  x8, x3, 2047
			32'h20 : Rom_data = 32'h00409493;	//slli  x9, x1, 4   
			32'h24 : Rom_data = 32'h0041d513;	//srli  x10, x3, 4
			32'h28 : Rom_data = 32'h4041d593;	//srai  x11, x3, 4
            default: Rom_data = 32'h00000013;   //NOP	
        endcase
    end
endmodule

